// Program memory implemented as combinational logic
// On the iCE40, this will be implemented in the logic fabric

// This is only used for the single-cycle machine; once we move to the
// multi-cycle design we will have a unified (and clocked) memory.

module progmem(input logic[31:0] addr,
               output logic[31:0] instr);

    // In the future, we will implement this by reading instructions stored in
    // an external file (which could be generated by an assembler), but for now
    // just hard-code the instructions here.
    // You can use Ripes to generate the bytes for the instructions you'd like
    // to run.

    always_comb
      case(addr)
        32'h0:  instr = 32'h00000013; // This is a NOP instruction (aka addi, x0, x0, 0)
        32'h4:  instr = 32'h001000b3; // Erase memory addy in x1 (aka addi x1, x0, x1)
        32'h8:  instr = 32'h00408093; // Adds 4 to register's self (addi x1, x1, 4)
        32'hc:  instr = 32'h00208133; // add x2 x1 x2 
        32'h10: instr = 32'h00108093; // Adds 1 to register's self (addi x1, x1, 1)
		32'h14: instr = 32'hfff08093; // addi x1 x1 -1
		32'h18: instr = 32'h001170b3; // and x1 x2 x1
		32'h1c: instr = 32'h001160b3; // or x1 x2 x1
		32'h20: instr = 32'h001140b3; // xor x1 x2 x1
		32'h24: instr = 32'h001120b3; //slt x1 x2 x1
		32'h28: instr = 32'h001130b3; // sltu x1 x2 x1
		32'h2c: instr = 32'h001110b3; // sll x1 x2 x1
		32'h30: instr = 32'h001150b3; // srl x1 x2 x1
		32'h34: instr = 32'h001100b3; // sub x1, x2, x1
		32'h38: instr = 32'h401150b3; // sra x1,x2,x1
      default: instr = 0;
    endcase

endmodule

